

***********************************
* TOP Circuit                     *
***********************************
.SUBCKT dco_model reset_ coarse_0  coarse_1  coarse_2  coarse_3  coarse_4  coarse_5  coarse_6  coarse_7  coarse_8  coarse_9   coarse_10  coarse_11  coarse_12  coarse_13  coarse_14  coarse_15  coarse_16  coarse_17  coarse_18  coarse_19   coarse_20  coarse_21  coarse_22  coarse_23  coarse_24  coarse_25  coarse_26  coarse_27  coarse_28  coarse_29   coarse_30  coarse_31  coarse_32  coarse_33  coarse_34  coarse_35  coarse_36  coarse_37  coarse_38  coarse_39   coarse_40  coarse_41  coarse_42  coarse_43  coarse_44  coarse_45  coarse_46  coarse_47  coarse_48  coarse_49   coarse_50  coarse_51  coarse_52  coarse_53  coarse_54  coarse_55  coarse_56  coarse_57  coarse_58  coarse_59   coarse_60  coarse_61  coarse_62  coarse_63  coarse_64  coarse_65  coarse_66  coarse_67  coarse_68  coarse_69   coarse_70  coarse_71  coarse_72  coarse_73  coarse_74  coarse_75  coarse_76  coarse_77  coarse_78  coarse_79   coarse_80  coarse_81  coarse_82  coarse_83  coarse_84  coarse_85  coarse_86  coarse_87  coarse_88  coarse_89   coarse_90  coarse_91  coarse_92  coarse_93  coarse_94  coarse_95  coarse_96  coarse_97  coarse_98  coarse_99   coarse_100  coarse_101  coarse_102  coarse_103  coarse_104  coarse_105  coarse_106  coarse_107  coarse_108  coarse_109   coarse_110  coarse_111  coarse_112  coarse_113  coarse_114  coarse_115  coarse_116  coarse_117  coarse_118  coarse_119   coarse_120  coarse_121  coarse_122  coarse_123  coarse_124  coarse_125  coarse_126  coarse_127  dco_out


XH000	reset_	dco_out	LINE1	AND2X1

XG000	coarse_0	LINE1	LINE2	TBUFIX4
XG001	coarse_1	LINE2	LINE3	TBUFIX4
XG002	coarse_2	LINE3	dco_out	TBUFIX4
XG003	coarse_3	LINE1	LINE2	TBUFIX4
XG004	coarse_4	LINE2	LINE3	TBUFIX4
XG005	coarse_5	LINE3	dco_out	TBUFIX4
XG006	coarse_6	LINE1	LINE2	TBUFIX4
XG007	coarse_7	LINE2	LINE3	TBUFIX4
XG008	coarse_8	LINE3	dco_out	TBUFIX4
XG009	coarse_9	LINE1	LINE2	TBUFIX4
XG010	coarse_10	LINE2	LINE3	TBUFIX4
XG011	coarse_11	LINE3	dco_out	TBUFIX4
XG012	coarse_12	LINE1	LINE2	TBUFIX4
XG013	coarse_13	LINE2	LINE3	TBUFIX4
XG014	coarse_14	LINE3	dco_out	TBUFIX4
XG015	coarse_15	LINE1	LINE2	TBUFIX4
XG016	coarse_16	LINE2	LINE3	TBUFIX4
XG017	coarse_17	LINE3	dco_out	TBUFIX4
XG018	coarse_18	LINE1	LINE2	TBUFIX4
XG019	coarse_19	LINE2	LINE3	TBUFIX4
XG020	coarse_20	LINE3	dco_out	TBUFIX4
XG021	coarse_21	LINE1	LINE2	TBUFIX4
XG022	coarse_22	LINE2	LINE3	TBUFIX4
XG023	coarse_23	LINE3	dco_out	TBUFIX4
XG024	coarse_24	LINE1	LINE2	TBUFIX4
XG025	coarse_25	LINE2	LINE3	TBUFIX4
XG026	coarse_26	LINE3	dco_out	TBUFIX4
XG027	coarse_27	LINE1	LINE2	TBUFIX4
XG028	coarse_28	LINE2	LINE3	TBUFIX4
XG029	coarse_29	LINE3	dco_out	TBUFIX4
XG030	coarse_30	LINE1	LINE2	TBUFIX4
XG031	coarse_31	LINE2	LINE3	TBUFIX4
XG032	coarse_32	LINE3	dco_out	TBUFIX4
XG033	coarse_33	LINE1	LINE2	TBUFIX4
XG034	coarse_34	LINE2	LINE3	TBUFIX4
XG035	coarse_35	LINE3	dco_out	TBUFIX4
XG036	coarse_36	LINE1	LINE2	TBUFIX4
XG037	coarse_37	LINE2	LINE3	TBUFIX4
XG038	coarse_38	LINE3	dco_out	TBUFIX4
XG039	coarse_39	LINE1	LINE2	TBUFIX4
XG040	coarse_40	LINE2	LINE3	TBUFIX4
XG041	coarse_41	LINE3	dco_out	TBUFIX4
XG042	coarse_42	LINE1	LINE2	TBUFIX4
XG043	coarse_43	LINE2	LINE3	TBUFIX4
XG044	coarse_44	LINE3	dco_out	TBUFIX4
XG045	coarse_45	LINE1	LINE2	TBUFIX4
XG046	coarse_46	LINE2	LINE3	TBUFIX4
XG047	coarse_47	LINE3	dco_out	TBUFIX4
XG048	coarse_48	LINE1	LINE2	TBUFIX4
XG049	coarse_49	LINE2	LINE3	TBUFIX4
XG050	coarse_50	LINE3	dco_out	TBUFIX4
XG051	coarse_51	LINE1	LINE2	TBUFIX4
XG052	coarse_52	LINE2	LINE3	TBUFIX4
XG053	coarse_53	LINE3	dco_out	TBUFIX4
XG054	coarse_54	LINE1	LINE2	TBUFIX4
XG055	coarse_55	LINE2	LINE3	TBUFIX4
XG056	coarse_56	LINE3	dco_out	TBUFIX4
XG057	coarse_57	LINE1	LINE2	TBUFIX4
XG058	coarse_58	LINE2	LINE3	TBUFIX4
XG059	coarse_59	LINE3	dco_out	TBUFIX4
XG060	coarse_60	LINE1	LINE2	TBUFIX4
XG061	coarse_61	LINE2	LINE3	TBUFIX4
XG062	coarse_62	LINE3	dco_out	TBUFIX4
XG063	coarse_63	LINE1	LINE2	TBUFIX4
XG064	coarse_64	LINE2	LINE3	TBUFIX4
XG065	coarse_65	LINE3	dco_out	TBUFIX4
XG066	coarse_66	LINE1	LINE2	TBUFIX4
XG067	coarse_67	LINE2	LINE2	TBUFIX4
XG068	coarse_68	LINE3	dco_out	TBUFIX4
XG069	coarse_69	LINE1	LINE2	TBUFIX4
XG070	coarse_70	LINE2	LINE3	TBUFIX4
XG071	coarse_71	LINE3	dco_out	TBUFIX4
XG072	coarse_72	LINE1	LINE2	TBUFIX4
XG073	coarse_73	LINE2	LINE3	TBUFIX4
XG074	coarse_74	LINE3	dco_out	TBUFIX4
XG075	coarse_75	LINE1	LINE2	TBUFIX4
XG076	coarse_76	LINE2	LINE3	TBUFIX4
XG077	coarse_77	LINE3	dco_out	TBUFIX4
XG078	coarse_78	LINE1	LINE2	TBUFIX4
XG079	coarse_79	LINE2	LINE3	TBUFIX4
XG080	coarse_80	LINE3	dco_out	TBUFIX4
XG081	coarse_81	LINE1	LINE2	TBUFIX4
XG082	coarse_82	LINE2	LINE3	TBUFIX4
XG083	coarse_83	LINE3	dco_out	TBUFIX4
XG084	coarse_84	LINE1	LINE2	TBUFIX4
XG085	coarse_85	LINE2	LINE3	TBUFIX4
XG086	coarse_86	LINE3	dco_out	TBUFIX4
XG087	coarse_87	LINE1	LINE2	TBUFIX4
XG088	coarse_88	LINE2	LINE3	TBUFIX4
XG089	coarse_89	LINE3	dco_out	TBUFIX4
XG090	coarse_90	LINE1	LINE2	TBUFIX4
XG091	coarse_91	LINE2	LINE3	TBUFIX4
XG092	coarse_92	LINE3	dco_out	TBUFIX4
XG093	coarse_93	LINE1	LINE2	TBUFIX4
XG094	coarse_94	LINE2	LINE3	TBUFIX4
XG095	coarse_95	LINE3	dco_out	TBUFIX4
XG096	coarse_96	LINE1	LINE2	TBUFIX4
XG097	coarse_97	LINE2	LINE3	TBUFIX4
XG098	coarse_98	LINE3	dco_out	TBUFIX4
XG099	coarse_99	LINE1	LINE2	TBUFIX4
XG100	coarse_100	LINE2	LINE3	TBUFIX4
XG101	coarse_101	LINE3	dco_out	TBUFIX4
XG102	coarse_102	LINE1	LINE2	TBUFIX4
XG103	coarse_103	LINE2	LINE3	TBUFIX4
XG104	coarse_104	LINE3	dco_out	TBUFIX4
XG105	coarse_105	LINE1	LINE2	TBUFIX4
XG106	coarse_106	LINE2	LINE3	TBUFIX4
XG107	coarse_107	LINE3	dco_out	TBUFIX4
XG108	coarse_108	LINE1	LINE2	TBUFIX4
XG109	coarse_109	LINE2	LINE3	TBUFIX4
XG110	coarse_110	LINE3	dco_out	TBUFIX4
XG111	coarse_111	LINE1	LINE2	TBUFIX4
XG112	coarse_112	LINE2	LINE3	TBUFIX4
XG113	coarse_113	LINE3	dco_out	TBUFIX4
XG114	coarse_114	LINE1	LINE2	TBUFIX4
XG115	coarse_115	LINE2	LINE3	TBUFIX4
XG116	coarse_116	LINE3	dco_out	TBUFIX4
XG117	coarse_117	LINE1	LINE2	TBUFIX4
XG118	coarse_118	LINE2	LINE3	TBUFIX4
XG119	coarse_119	LINE3	dco_out	TBUFIX4
XG120	coarse_120	LINE1	LINE2	TBUFIX4
XG121	coarse_121	LINE2	LINE3	TBUFIX4
XG122	coarse_122	LINE3	dco_out	TBUFIX4
XG123	coarse_123	LINE1	LINE2	TBUFIX4
XG124	coarse_124	LINE2	LINE3	TBUFIX4
XG125	coarse_125	LINE3	dco_out	TBUFIX4
XG126	coarse_126	LINE1	LINE2	TBUFIX4
XG127	coarse_127	LINE2	LINE2	TBUFIX4



C1    dco_out    0 0.02p
.ENDS 
***********************************
* Subckt Definition               *
***********************************
.SUBCKT INVERTER Y A pl=0.24u pw=0.24u nl=0.24u nw=0.24u
M_N   Y  A VSS VSS N_18_G2 w=nw l=nl
M_P VDD  A   Y VDD P_18_G2 w=pw l=pl
.ENDS INVERTER

.end
